package piso_types;
parameter int timeout_delay_p = 8;
parameter int pbytes_p = 4;
parameter int pwidth_p = pbytes_p * 8;

typedef logic [1:0] pbyte_count_t;


endpackage : piso_types
